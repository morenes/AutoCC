bind dcp_pipe dcp_pipe_prop
	#(
		.ASSERT_INPUTS (0)
	) u_dcp_pipe_sva(.*);