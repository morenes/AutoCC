bind is_core_wrap is_core_prop
	#(
		.ASSERT_INPUTS (0)
	) u_is_core_sva(.*);