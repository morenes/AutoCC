bind cva6_wrap cva6_prop
	#(
		.ASSERT_INPUTS (0)
	) u_cva6_sva(.*);